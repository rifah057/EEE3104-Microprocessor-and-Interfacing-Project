module tb_full();
  reg clk;
  reg reset;
  wire Cp, Ep, Lmp, Lmi, Cei, Cea, Li, Ei, LaRam, Lab, LaALU, Eatmp, Lbtmp, Ltmpa, Etmpb, Su, Eu, Eba, Lo, EaRAM, LA, LtmpRAM, Cetmp, LbALU, LaOUT, EaOut;
  wire[3:0] PC_to_MAR; // connection between pc to mar
  wire[3:0] MAR_to_RAM; //connection between mar to ram
  wire[7:0] RAM_to_IR; //connection between ram and ir
  wire[3:0] RAM_to_A; //connection between ram and a
  wire[3:0] IR_to_Control; //connection between ir and control unit
  wire[3:0] IR_to_MAR; //connection between ir and mar
  wire[3:0] A_to_ALU; //connection between a and alu
  wire[3:0] B_to_A; //connection between a and b
  wire[3:0] A_to_TMP; //connection between a and temp
  wire[3:0] TMP_to_B; //connection between tmp and b
  wire[3:0] B_to_ALU; //connection between b and alu
  wire[3:0] ALU_to_A; //connection between a and alu
  wire[3:0] A_to_RAM; //connection between a and ram(to send data to ram from A)
  wire[3:0] RAM_to_TMP; //connection between ram and tmp
  wire[3:0] ALU_to_B; //connection between alu and b(to send data from alu to b)
  wire[3:0] TMP_to_ALU; //connection between tmp and alu
  wire[3:0] A_to_OUT; //connection between a and out
  wire[3:0] OUT_to_disp; //connection between out and display
  
  ControlSequencer example_tbCS(clk, reset, IR_to_Control, Cp, Ep, Lmp, Lmi, Cei, Cea, Li, Ei, LaRam, Lab, LaALU, Eatmp, Su, Eu, Lbtmp, Eba, Lo, Ltmpa, Etmpb, EaRAM, LA, LtmpRAM, Cetmp, LbALU, LaOUT, EaOut);
  ProgramCounter example_tbPC(clk, reset, Ep, Cp, PC_to_MAR);
  MAR example_tbMAR(clk, Lmp, Lmi, PC_to_MAR, IR_to_MAR, MAR_to_RAM);
  RAM example_tbRAMRAM(clk, Cei, Cea, Cetmp, LA, MAR_to_RAM, RAM_to_IR, RAM_to_A, A_to_RAM, RAM_to_A);
  InstructionRegister example_tbIR(clk, RAM_to_IR, Li, Ei, reset, IR_to_Control, IR_to_MAR);
  ARegister example_tbAR(clk, RAM_to_A, B_to_A, LaRam, Lab, LaALU, Eatmp, EaRAM, EaOut, reset, A_to_ALU, A_to_TMP, ALU_to_A, A_to_RAM, A_to_OUT);
  TMPRegister example_tbTMPR(clk, A_to_TMP, Ltmpa, LtmpRAM, Etmpb, reset, TMP_to_B, RAM_to_TMP);
  BRegister example_tbBR(clk, TMP_to_B, Lbtmp, LbALU, Eba, reset, B_to_A, B_to_ALU, ALU_to_B);
  ALU example_tbALU(clk, reset, A_to_ALU, B_to_ALU, TMP_to_ALU, IR_to_Control, Eu, ALU_to_A, ALU_to_B);
  OUTRegister example_tbOUTR(clk, reset, A_to_OUT, LaOUT, OUT_to_disp);

  initial
    begin
      clk = 1'b1;
      reset = 1'b1; 
      #1 reset = 1'b0; //reset is done once
      #2 $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #1 reset = 1'b1;
      #3
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A);
      
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM);
      
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM);
      
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM);
      
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM);
      
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM);
      
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM);
      
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM);
      
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM);
      
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, LtmpRAM=%b, Cetmp=%b, LbALU=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b, RAM_to_TMP=%4b, TMP_to_ALU=%4b, ALU_to_B=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, LtmpRAM, Cetmp, LbALU, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM, RAM_to_TMP, TMP_to_ALU, ALU_to_B);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, LtmpRAM=%b, Cetmp=%b, LbALU=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b, RAM_to_TMP=%4b, TMP_to_ALU=%4b, ALU_to_B=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, LtmpRAM, Cetmp, LbALU, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM, RAM_to_TMP, TMP_to_ALU, ALU_to_B);
      
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, LtmpRAM=%b, Cetmp=%b, LbALU=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b, RAM_to_TMP=%4b, TMP_to_ALU=%4b, ALU_to_B=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, LtmpRAM, Cetmp, LbALU, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM, RAM_to_TMP, TMP_to_ALU, ALU_to_B);
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, LtmpRAM=%b, Cetmp=%b, LbALU=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b, RAM_to_TMP=%4b, TMP_to_ALU=%4b, ALU_to_B=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, LtmpRAM, Cetmp, LbALU, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM, RAM_to_TMP, TMP_to_ALU, ALU_to_B);
      
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, LtmpRAM=%b, Cetmp=%b, LbALU=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b, RAM_to_TMP=%4b, TMP_to_ALU=%4b, ALU_to_B=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, LtmpRAM, Cetmp, LbALU, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM, RAM_to_TMP, TMP_to_ALU, ALU_to_B);
      
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, LtmpRAM=%b, Cetmp=%b, LbALU=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b, RAM_to_TMP=%4b, TMP_to_ALU=%4b, ALU_to_B=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, LtmpRAM, Cetmp, LbALU, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM, RAM_to_TMP, TMP_to_ALU, ALU_to_B);
      
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, LtmpRAM=%b, Cetmp=%b, LbALU=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b, RAM_to_TMP=%4b, TMP_to_ALU=%4b, ALU_to_B=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, LtmpRAM, Cetmp, LbALU, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM, RAM_to_TMP, TMP_to_ALU, ALU_to_B);
      
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, LtmpRAM=%b, Cetmp=%b, LbALU=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b, RAM_to_TMP=%4b, TMP_to_ALU=%4b, ALU_to_B=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, LtmpRAM, Cetmp, LbALU, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM, RAM_to_TMP, TMP_to_ALU, ALU_to_B);
      
      
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, LtmpRAM=%b, Cetmp=%b, LbALU=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b, RAM_to_TMP=%4b, TMP_to_ALU=%4b, ALU_to_B=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, LtmpRAM, Cetmp, LbALU, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM, RAM_to_TMP, TMP_to_ALU, ALU_to_B);
      
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, LtmpRAM=%b, Cetmp=%b, LbALU=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b, RAM_to_TMP=%4b, TMP_to_ALU=%4b, ALU_to_B=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, LtmpRAM, Cetmp, LbALU, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM, RAM_to_TMP, TMP_to_ALU, ALU_to_B);
      
      
      
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, LtmpRAM=%b, Cetmp=%b, LbALU=%b, LaOUT=%b, EaOut=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b, RAM_to_TMP=%4b, TMP_to_ALU=%4b, ALU_to_B=%4b, A_to_OUT=%4b, OUT_to_disp=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, LtmpRAM, Cetmp, LbALU, LaOUT, EaOut, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM, RAM_to_TMP, TMP_to_ALU, ALU_to_B, A_to_OUT, OUT_to_disp);
      
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, LtmpRAM=%b, Cetmp=%b, LbALU=%b, LaOUT=%b, EaOut=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b, RAM_to_TMP=%4b, TMP_to_ALU=%4b, ALU_to_B=%4b, A_to_OUT=%4b, OUT_to_disp=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, LtmpRAM, Cetmp, LbALU, LaOUT, EaOut, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM, RAM_to_TMP, TMP_to_ALU, ALU_to_B, A_to_OUT, OUT_to_disp);
      
      #4
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, LtmpRAM=%b, Cetmp=%b, LbALU=%b, LaOUT=%b, EaOut=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b, RAM_to_TMP=%4b, TMP_to_ALU=%4b, ALU_to_B=%4b, A_to_OUT=%4b, OUT_to_disp=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, LtmpRAM, Cetmp, LbALU, LaOUT, EaOut, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM, RAM_to_TMP, TMP_to_ALU, ALU_to_B, A_to_OUT, OUT_to_disp);
      
      #6
      $display("t=%d, Cp=%b, Ep=%b, Cei=%b, Cea=%b, LaRam=%b, Lab=%b, Eba=%b, Eatmp=%b, Lbtmp=%b, Ltmpa=%b, Etmpb=%b, Ei=%b, Li=%b, Lmp = %b, Lmi=%b, Su=%b, LaALU=%4b, Eu=%b, Lo=%b, LA=%b, EaRAM=%b, LtmpRAM=%b, Cetmp=%b, LbALU=%b, LaOUT=%b, EaOut=%b, PC_to_MAR=%8b, MAR_to_RAM=%8b, RAM_to_IR=%8b, IR_to_Control=%4b, IR_to_MAR=%4b, RAM_to_A=%4b, A_to_ALU=%4b, A_to_TMP=%4b, TMP_to_B=%4b, B_to_A=%4b, ALU_to_A=%4b, A_to_RAM=%4b, RAM_to_TMP=%4b, TMP_to_ALU=%4b, ALU_to_B=%4b, A_to_OUT=%4b, OUT_to_disp=%4b", $time, Cp, Ep, Cei, Cea, LaRam, Lab, Eba, Eatmp, Lbtmp, Ltmpa, Etmpb, Ei, Li, Lmp, Lmi, Su, LaALU, Eu, Lo, LA, EaRAM, LtmpRAM, Cetmp, LbALU, LaOUT, EaOut, PC_to_MAR, MAR_to_RAM, RAM_to_IR, IR_to_Control, IR_to_MAR, RAM_to_A, A_to_ALU, A_to_TMP, TMP_to_B, B_to_A, ALU_to_A, A_to_RAM, RAM_to_TMP, TMP_to_ALU, ALU_to_B, A_to_OUT, OUT_to_disp);
      
      
      #5
      $finish;
    end
  
  always #5 clk = ~clk;

endmodule    

